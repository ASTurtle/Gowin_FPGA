module testfft_top (
    input clk,
    input reset_n,
    output [55:1] out,
    input  [40:1] in
);





endmodule