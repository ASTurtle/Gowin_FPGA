`define MODULE_NAME Equalizer
`define MUL_5;
